// Code your design here
module notgate(Y,A);
  input A;
  output Y;
  assign Y=~A;
endmodule
